Library ieee;
use ieee.std_logic_1164.all;

entity serrure_Tb is

end serrure_Tb ;

architecture arc_serrure_Tb of serrure_Tb is

signal ch1,ch2,ch3,ch4 : std_logic_vector(15 downto 0);
signal clock :  std_logic ;
signal clear :  std_logic ;
signal writ : std_logic ;
signal S1,S2,S3,S4 :  std_logic_vector(3 downto 0);
signal S5,S6,S7,S8 : std_logic; 
signal s : std_logic_vector(15 downto 0);
signal r : std_logic ;

component serrure 
port(
    chiffre1 : in std_logic_vector(15 downto 0);
    chiffre2 : in std_logic_vector(15 downto 0);
    chiffre3 : in std_logic_vector(15 downto 0);
    chiffre4 : in std_logic_vector(15 downto 0);
    w : in std_logic ;
    clock : in std_logic ;
    clear : in std_logic ;
    sortie : out std_logic_vector(15 downto 0);
    Sb1,Sb2,Sb3,Sb4 : out std_logic_vector(3 downto 0);
    Sb5,Sb6,Sb7,Sb8 : out std_logic ;
    S : out std_logic 
);
end component ;

begin
inst : serrure port map(ch1,ch2,ch3,ch4,writ,clock,clear,s,S1,S2,S3,S4,S5,S6,S7,S8,r);
process
begin
ch1 <= "0000000000000000";
ch2 <= "0000000000000000";
ch3 <= "0000000000000000";
ch4 <= "0000000000000000";
wait for 20 ns;
ch1 <= "0000000000000001";
ch2 <= "0000000000000010";
ch3 <= "0000000000000100";
ch4 <= "0000000000010000";
wait for 300 ns;
ch1 <= "0000000000000000";
ch2 <= "0000000000000000";
ch3 <= "0000000000000000";
ch4 <= "0000000000000000";
wait for 100 ns;
ch1 <= "0000000000100000";
ch2 <= "0000000001000000";
ch3 <= "0000000100000000";
ch4 <= "0000001000000000";
wait for 300 ns;
ch1 <= "0000000000000000";
ch2 <= "0000000000000000";
ch3 <= "0000000000000000";
ch4 <= "0000000000000000";
wait for 100 ns;
ch1 <= "0000000000000001";
ch2 <= "0000000000000010";
ch3 <= "0000000000000100";
ch4 <= "0000000000010000";
wait for 300 ns;
ch1 <= "0000000000000000";
ch2 <= "0000000000000000";
ch3 <= "0000000000000000";
ch4 <= "0000000000000000";
wait;

end process;

process
begin
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait for 10 ns;
clock <= '1';
wait for 10 ns;
clock <= '0';
wait;
end process;

process

begin
clear <= '1';
wait for 110 ns;
clear <= '0';
wait for 200 ns;
clear <= '1';
wait for 200 ns;
clear <= '0';
wait for 200 ns;
clear <= '1';
wait for 200 ns;
clear <= '0';
wait for 200 ns;
clear <= '1';
wait for 200 ns;
clear <= '0';
wait for 200 ns;
clear <= '1';
wait for 200 ns;
clear <= '0';
wait for 200 ns;
clear <= '1';
wait for 200 ns;
clear <= '0';
wait for 200 ns;
clear <= '1';
wait for 200 ns;
clear <= '0';
wait for 200 ns;
clear <= '1';
wait;

end process;

process 
begin
writ <= '1';
wait ;
end process;

end arc_serrure_Tb;
